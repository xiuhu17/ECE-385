module control (	);
						
	   
	
endmodule