module S_BOX_MAP(input logic[47:0] input_data,
                 output logic[31:0] output_data);
    parameter [3:0]S_BOX_ROM[8][4][16] = {
        {
            {{14},{4},{13},{1},{2},{15},{11},{8},{3},{10},{6},{12},{5},{9},{0},{7}},
            {{0},{15},{7},{4},{14},{2},{13},{1},{10},{6},{12},{11},{9},{5},{3},{8}},
            {{4},{1},{14},{8},{13},{6},{2},{11},{15},{12},{9},{7},{3},{10},{5},{0}},
            {{15},{12},{8},{2},{4},{9},{1},{7},{5},{11},{3},{14},{10},{0},{6},{13}}
        },
        {
            {{15},{1},{8},{14},{6},{11},{3},{4},{9},{7},{2},{13},{12},{0},{5},{10}},
            {{3},{13},{4},{7},{15},{2},{8},{14},{12},{0},{1},{10},{6},{9},{11},{5}},
            {{0},{14},{7},{11},{10},{4},{13},{1},{5},{8},{12},{6},{9},{3},{2},{15}},
            {{13},{8},{10},{1},{3},{15},{4},{2},{11},{6},{7},{12},{0},{5},{14},{9}}
        },
        {
            {{10},{0},{9},{14},{6},{3},{15},{5},{1},{13},{12},{7},{11},{4},{2},{8}},
            {{13},{7},{0},{9},{3},{4},{6},{10},{2},{8},{5},{14},{12},{11},{15},{1}},
            {{13},{6},{4},{9},{8},{15},{3},{0},{11},{1},{2},{12},{5},{10},{14},{7}},
            {{1},{10},{13},{0},{6},{9},{8},{7},{4},{15},{14},{3},{11},{5},{2},{12}}
        },
        {
            {{7},{13},{14},{3},{0},{6},{9},{10},{1},{2},{8},{5},{11},{12},{4},{15}},
            {{13},{8},{11},{5},{6},{15},{0},{3},{4},{7},{2},{12},{1},{10},{14},{9}},
            {{10},{6},{9},{0},{12},{11},{7},{13},{15},{1},{3},{14},{5},{2},{8},{4}},
            {{3},{15},{0},{6},{10},{1},{13},{8},{9},{4},{5},{11},{12},{7},{2},{14}}
        },
        {
            {{2},{12},{4},{1},{7},{10},{11},{6},{8},{5},{3},{15},{13},{0},{14},{9}},
            {{14},{11},{2},{12},{4},{7},{13},{1},{5},{0},{15},{10},{3},{9},{8},{6}},
            {{4},{2},{1},{11},{10},{13},{7},{8},{15},{9},{12},{5},{6},{3},{0},{14}},
            {{11},{8},{12},{7},{1},{14},{2},{13},{6},{15},{0},{9},{10},{4},{5},{3}}
        },
        {
            {{12},{1},{10},{15},{9},{2},{6},{8},{0},{13},{3},{4},{14},{7},{5},{11}},
            {{10},{15},{4},{2},{7},{12},{9},{5},{6},{1},{13},{14},{0},{11},{3},{8}},
            {{9},{14},{15},{5},{2},{8},{12},{3},{7},{0},{4},{10},{1},{13},{11},{6}},
            {{4},{3},{2},{12},{9},{5},{15},{10},{11},{14},{1},{7},{6},{0},{8},{13}}
        },
        {
            {{4},{11},{2},{14},{15},{0},{8},{13},{3},{12},{9},{7},{5},{10},{6},{1}},
            {{13},{0},{11},{7},{4},{9},{1},{10},{14},{3},{5},{12},{2},{15},{8},{6}},
            {{1},{4},{11},{13},{12},{3},{7},{14},{10},{15},{6},{8},{0},{5},{9},{2}},
            {{6},{11},{13},{8},{1},{4},{10},{7},{9},{5},{0},{15},{14},{2},{3},{12}}
        },
        
        {
            {{13},{2},{8},{4},{6},{15},{11},{1},{10},{9},{3},{14},{5},{0},{12},{7}},
            {{1},{15},{13},{8},{10},{3},{7},{4},{12},{5},{6},{11},{0},{14},{9},{2}},
            {{7},{11},{4},{1},{9},{12},{14},{2},{0},{6},{10},{13},{15},{3},{5},{8}},
            {{2},{1},{14},{7},{4},{10},{8},{13},{15},{12},{9},{0},{3},{5},{6},{11}}
        }
    };

    logic [1:0] row0, row1, row2, row3, row4, row5, row6, row7;
    assign row0 = {{input_data[47]}, {input_data[42]}};
    assign row1 = {{input_data[41]}, {input_data[36]}};
    assign row2 = {{input_data[35]}, {input_data[30]}};
    assign row3 = {{input_data[29]}, {input_data[24]}};
    assign row4 = {{input_data[23]}, {input_data[18]}};
    assign row5 = {{input_data[17]}, {input_data[12]}};
    assign row6 = {{input_data[11]}, {input_data[6]}};
    assign row7 = {{input_data[5]}, {input_data[0]}};


    assign output_data = {
        {S_BOX_ROM[row0][input_data[46:43]]},
        {S_BOX_ROM[row1][input_data[40:37]]},
        {S_BOX_ROM[row2][input_data[34:31]]},
        {S_BOX_ROM[row3][input_data[28:25]]},
        {S_BOX_ROM[row4][input_data[22:19]]},
        {S_BOX_ROM[row5][input_data[16:13]]},
        {S_BOX_ROM[row6][input_data[10:7]]},
        {S_BOX_ROM[row7][input_data[4:1]]}
    };

endmodule