module P_BOX_Permutate();

endmodule