module CNTRL(output logic [3:0] red, green, blue);

endmodule